module charactermap (
           input wire clk,
           input wire [7:0] character,
           output reg [127:0] characterraster
       );

always @(posedge clk)
begin
    case (character)
        8'h00 : characterraster = 128'h00000000000000000000000000000000;
        8'h01 : characterraster = 128'h00007E81A58181BD9981817E00000000;
        8'h02 : characterraster = 128'h00007EFFDBFFFFC3E7FFFF7E00000000;
        8'h03 : characterraster = 128'h000000006CFEFEFEFE7C381000000000;
        8'h04 : characterraster = 128'h0000000010387CFE7C38100000000000;
        8'h05 : characterraster = 128'h000000183C3CE7E7E718183C00000000;
        8'h06 : characterraster = 128'h000000183C7EFFFF7E18183C00000000;
        8'h07 : characterraster = 128'h000000000000183C3C18000000000000;
        8'h08 : characterraster = 128'hFFFFFFFFFFFFE7C3C3E7FFFFFFFFFFFF;
        8'h09 : characterraster = 128'h00000000003C664242663C0000000000;
        8'h0A : characterraster = 128'hFFFFFFFFFFC399BDBD99C3FFFFFFFFFF;
        8'h0B : characterraster = 128'h00001E0E1A3278CCCCCCCC7800000000;
        8'h0C : characterraster = 128'h00003C666666663C187E181800000000;
        8'h0D : characterraster = 128'h00003F333F3030303070F0E000000000;
        8'h0E : characterraster = 128'h00007F637F6363636367E7E6C0000000;
        8'h0F : characterraster = 128'h0000001818DB3CE73CDB181800000000;
        8'h10 : characterraster = 128'h0080C0E0F0F8FEF8F0E0C08000000000;
        8'h11 : characterraster = 128'h0002060E1E3EFE3E1E0E060200000000;
        8'h12 : characterraster = 128'h0000183C7E1818187E3C180000000000;
        8'h13 : characterraster = 128'h00006666666666666600666600000000;
        8'h14 : characterraster = 128'h00007FDBDBDB7B1B1B1B1B1B00000000;
        8'h15 : characterraster = 128'h007CC660386CC6C66C380CC67C000000;
        8'h16 : characterraster = 128'h0000000000000000FEFEFEFE00000000;
        8'h17 : characterraster = 128'h0000183C7E1818187E3C187E00000000;
        8'h18 : characterraster = 128'h0000183C7E1818181818181800000000;
        8'h19 : characterraster = 128'h0000181818181818187E3C1800000000;
        8'h1A : characterraster = 128'h0000000000180CFE0C18000000000000;
        8'h1B : characterraster = 128'h00000000003060FE6030000000000000;
        8'h1C : characterraster = 128'h000000000000C0C0C0FE000000000000;
        8'h1D : characterraster = 128'h0000000000286CFE6C28000000000000;
        8'h1E : characterraster = 128'h000000001038387C7CFEFE0000000000;
        8'h1F : characterraster = 128'h00000000FEFE7C7C3838100000000000;
        8'h20 : characterraster = 128'h00000000000000000000000000000000;
        8'h21 : characterraster = 128'h0000183C3C3C18181800181800000000;
        8'h22 : characterraster = 128'h00666666240000000000000000000000;
        8'h23 : characterraster = 128'h0000006C6CFE6C6C6CFE6C6C00000000;
        8'h24 : characterraster = 128'h18187CC6C2C07C060686C67C18180000;
        8'h25 : characterraster = 128'h00000000C2C60C183060C68600000000;
        8'h26 : characterraster = 128'h0000386C6C3876DCCCCCCC7600000000;
        8'h27 : characterraster = 128'h00303030600000000000000000000000;
        8'h28 : characterraster = 128'h00000C18303030303030180C00000000;
        8'h29 : characterraster = 128'h000030180C0C0C0C0C0C183000000000;
        8'h2A : characterraster = 128'h0000000000663CFF3C66000000000000;
        8'h2B : characterraster = 128'h000000000018187E1818000000000000;
        8'h2C : characterraster = 128'h00000000000000000018181830000000;
        8'h2D : characterraster = 128'h00000000000000FE0000000000000000;
        8'h2E : characterraster = 128'h00000000000000000000181800000000;
        8'h2F : characterraster = 128'h0000000002060C183060C08000000000;
        8'h30 : characterraster = 128'h0000386CC6C6D6D6C6C66C3800000000;
        8'h31 : characterraster = 128'h00001838781818181818187E00000000;
        8'h32 : characterraster = 128'h00007CC6060C183060C0C6FE00000000;
        8'h33 : characterraster = 128'h00007CC606063C060606C67C00000000;
        8'h34 : characterraster = 128'h00000C1C3C6CCCFE0C0C0C1E00000000;
        8'h35 : characterraster = 128'h0000FEC0C0C0FC060606C67C00000000;
        8'h36 : characterraster = 128'h00003860C0C0FCC6C6C6C67C00000000;
        8'h37 : characterraster = 128'h0000FEC606060C183030303000000000;
        8'h38 : characterraster = 128'h00007CC6C6C67CC6C6C6C67C00000000;
        8'h39 : characterraster = 128'h00007CC6C6C67E0606060C7800000000;
        8'h3A : characterraster = 128'h00000000181800000018180000000000;
        8'h3B : characterraster = 128'h00000000181800000018183000000000;
        8'h3C : characterraster = 128'h000000060C18306030180C0600000000;
        8'h3D : characterraster = 128'h00000000007E00007E00000000000000;
        8'h3E : characterraster = 128'h0000006030180C060C18306000000000;
        8'h3F : characterraster = 128'h00007CC6C60C18181800181800000000;
        8'h40 : characterraster = 128'h0000007CC6C6DEDEDEDCC07C00000000;
        8'h41 : characterraster = 128'h000010386CC6C6FEC6C6C6C600000000;
        8'h42 : characterraster = 128'h0000FC6666667C66666666FC00000000;
        8'h43 : characterraster = 128'h00003C66C2C0C0C0C0C2663C00000000;
        8'h44 : characterraster = 128'h0000F86C6666666666666CF800000000;
        8'h45 : characterraster = 128'h0000FE6662687868606266FE00000000;
        8'h46 : characterraster = 128'h0000FE6662687868606060F000000000;
        8'h47 : characterraster = 128'h00003C66C2C0C0DEC6C6663A00000000;
        8'h48 : characterraster = 128'h0000C6C6C6C6FEC6C6C6C6C600000000;
        8'h49 : characterraster = 128'h00003C18181818181818183C00000000;
        8'h4A : characterraster = 128'h00001E0C0C0C0C0CCCCCCC7800000000;
        8'h4B : characterraster = 128'h0000E666666C78786C6666E600000000;
        8'h4C : characterraster = 128'h0000F06060606060606266FE00000000;
        8'h4D : characterraster = 128'h0000C6EEFEFED6C6C6C6C6C600000000;
        8'h4E : characterraster = 128'h0000C6E6F6FEDECEC6C6C6C600000000;
        8'h4F : characterraster = 128'h00007CC6C6C6C6C6C6C6C67C00000000;
        8'h50 : characterraster = 128'h0000FC6666667C60606060F000000000;
        8'h51 : characterraster = 128'h00007CC6C6C6C6C6C6D6DE7C0C0E0000;
        8'h52 : characterraster = 128'h0000FC6666667C6C666666E600000000;
        8'h53 : characterraster = 128'h00007CC6C660380C06C6C67C00000000;
        8'h54 : characterraster = 128'h00007E7E5A1818181818183C00000000;
        8'h55 : characterraster = 128'h0000C6C6C6C6C6C6C6C6C67C00000000;
        8'h56 : characterraster = 128'h0000C6C6C6C6C6C6C66C381000000000;
        8'h57 : characterraster = 128'h0000C6C6C6C6D6D6D6FEEE6C00000000;
        8'h58 : characterraster = 128'h0000C6C66C7C38387C6CC6C600000000;
        8'h59 : characterraster = 128'h0000666666663C181818183C00000000;
        8'h5A : characterraster = 128'h0000FEC6860C183060C2C6FE00000000;
        8'h5B : characterraster = 128'h00003C30303030303030303C00000000;
        8'h5C : characterraster = 128'h00000080C0E070381C0E060200000000;
        8'h5D : characterraster = 128'h00003C0C0C0C0C0C0C0C0C3C00000000;
        8'h5E : characterraster = 128'h10386CC6000000000000000000000000;
        8'h5F : characterraster = 128'h00000000000000000000000000FF0000;
        8'h60 : characterraster = 128'h30301800000000000000000000000000;
        8'h61 : characterraster = 128'h0000000000780C7CCCCCCC7600000000;
        8'h62 : characterraster = 128'h0000E06060786C666666667C00000000;
        8'h63 : characterraster = 128'h00000000007CC6C0C0C0C67C00000000;
        8'h64 : characterraster = 128'h00001C0C0C3C6CCCCCCCCC7600000000;
        8'h65 : characterraster = 128'h00000000007CC6FEC0C0C67C00000000;
        8'h66 : characterraster = 128'h0000386C6460F060606060F000000000;
        8'h67 : characterraster = 128'h000000000076CCCCCCCCCC7C0CCC7800;
        8'h68 : characterraster = 128'h0000E060606C7666666666E600000000;
        8'h69 : characterraster = 128'h00001818003818181818183C00000000;
        8'h6A : characterraster = 128'h00000606000E06060606060666663C00;
        8'h6B : characterraster = 128'h0000E06060666C78786C66E600000000;
        8'h6C : characterraster = 128'h00003818181818181818183C00000000;
        8'h6D : characterraster = 128'h0000000000ECFED6D6D6D6C600000000;
        8'h6E : characterraster = 128'h0000000000DC66666666666600000000;
        8'h6F : characterraster = 128'h00000000007CC6C6C6C6C67C00000000;
        8'h70 : characterraster = 128'h0000000000DC66666666667C6060F000;
        8'h71 : characterraster = 128'h000000000076CCCCCCCCCC7C0C0C1E00;
        8'h72 : characterraster = 128'h0000000000DC7666606060F000000000;
        8'h73 : characterraster = 128'h00000000007CC660380CC67C00000000;
        8'h74 : characterraster = 128'h0000103030FC30303030361C00000000;
        8'h75 : characterraster = 128'h0000000000CCCCCCCCCCCC7600000000;
        8'h76 : characterraster = 128'h000000000066666666663C1800000000;
        8'h77 : characterraster = 128'h0000000000C6C6D6D6D6FE6C00000000;
        8'h78 : characterraster = 128'h0000000000C66C3838386CC600000000;
        8'h79 : characterraster = 128'h0000000000C6C6C6C6C6C67E060CF800;
        8'h7A : characterraster = 128'h0000000000FECC183060C6FE00000000;
        8'h7B : characterraster = 128'h00000E18181870181818180E00000000;
        8'h7C : characterraster = 128'h00001818181800181818181800000000;
        8'h7D : characterraster = 128'h0000701818180E181818187000000000;
        8'h7E : characterraster = 128'h000076DC000000000000000000000000;
        8'h7F : characterraster = 128'h0000000010386CC6C6C6FE0000000000;
        8'h80 : characterraster = 128'h00003C66C2C0C0C0C2663C0C067C0000;
        8'h81 : characterraster = 128'h0000CC0000CCCCCCCCCCCC7600000000;
        8'h82 : characterraster = 128'h000C1830007CC6FEC0C0C67C00000000;
        8'h83 : characterraster = 128'h0010386C00780C7CCCCCCC7600000000;
        8'h84 : characterraster = 128'h0000CC0000780C7CCCCCCC7600000000;
        8'h85 : characterraster = 128'h0060301800780C7CCCCCCC7600000000;
        8'h86 : characterraster = 128'h00386C3800780C7CCCCCCC7600000000;
        8'h87 : characterraster = 128'h000000003C666060663C0C063C000000;
        8'h88 : characterraster = 128'h0010386C007CC6FEC0C0C67C00000000;
        8'h89 : characterraster = 128'h0000C600007CC6FEC0C0C67C00000000;
        8'h8A : characterraster = 128'h00603018007CC6FEC0C0C67C00000000;
        8'h8B : characterraster = 128'h00006600003818181818183C00000000;
        8'h8C : characterraster = 128'h00183C66003818181818183C00000000;
        8'h8D : characterraster = 128'h00603018003818181818183C00000000;
        8'h8E : characterraster = 128'h00C60010386CC6C6FEC6C6C600000000;
        8'h8F : characterraster = 128'h386C3800386CC6C6FEC6C6C600000000;
        8'h90 : characterraster = 128'h18306000FE66607C606066FE00000000;
        8'h91 : characterraster = 128'h0000000000CC76367ED8D86E00000000;
        8'h92 : characterraster = 128'h00003E6CCCCCFECCCCCCCCCE00000000;
        8'h93 : characterraster = 128'h0010386C007CC6C6C6C6C67C00000000;
        8'h94 : characterraster = 128'h0000C600007CC6C6C6C6C67C00000000;
        8'h95 : characterraster = 128'h00603018007CC6C6C6C6C67C00000000;
        8'h96 : characterraster = 128'h003078CC00CCCCCCCCCCCC7600000000;
        8'h97 : characterraster = 128'h0060301800CCCCCCCCCCCC7600000000;
        8'h98 : characterraster = 128'h0000C60000C6C6C6C6C6C67E060C7800;
        8'h99 : characterraster = 128'h00C6007CC6C6C6C6C6C6C67C00000000;
        8'h9A : characterraster = 128'h00C600C6C6C6C6C6C6C6C67C00000000;
        8'h9B : characterraster = 128'h0018183C66606060663C181800000000;
        8'h9C : characterraster = 128'h00386C6460F060606060E6FC00000000;
        8'h9D : characterraster = 128'h000066663C187E187E18181800000000;
        8'h9E : characterraster = 128'h00F8CCCCF8C4CCDECCCCCCC600000000;
        8'h9F : characterraster = 128'h000E1B1818187E1818181818D8700000;
        8'hA0 : characterraster = 128'h0018306000780C7CCCCCCC7600000000;
        8'hA1 : characterraster = 128'h000C1830003818181818183C00000000;
        8'hA2 : characterraster = 128'h00183060007CC6C6C6C6C67C00000000;
        8'hA3 : characterraster = 128'h0018306000CCCCCCCCCCCC7600000000;
        8'hA4 : characterraster = 128'h000076DC00DC66666666666600000000;
        8'hA5 : characterraster = 128'h76DC00C6E6F6FEDECEC6C6C600000000;
        8'hA6 : characterraster = 128'h003C6C6C3E007E000000000000000000;
        8'hA7 : characterraster = 128'h00386C6C38007C000000000000000000;
        8'hA8 : characterraster = 128'h0000303000303060C0C6C67C00000000;
        8'hA9 : characterraster = 128'h000000000000FEC0C0C0C00000000000;
        8'hAA : characterraster = 128'h000000000000FE060606060000000000;
        8'hAB : characterraster = 128'h00C0C0C2C6CC183060DC860C183E0000;
        8'hAC : characterraster = 128'h00C0C0C2C6CC183066CE9E3E06060000;
        8'hAD : characterraster = 128'h00001818001818183C3C3C1800000000;
        8'hAE : characterraster = 128'h0000000000366CD86C36000000000000;
        8'hAF : characterraster = 128'h0000000000D86C366CD8000000000000;
        8'hB0 : characterraster = 128'h11441144114411441144114411441144;
        8'hB1 : characterraster = 128'h55AA55AA55AA55AA55AA55AA55AA55AA;
        8'hB2 : characterraster = 128'hDD77DD77DD77DD77DD77DD77DD77DD77;
        8'hB3 : characterraster = 128'h18181818181818181818181818181818;
        8'hB4 : characterraster = 128'h18181818181818F81818181818181818;
        8'hB5 : characterraster = 128'h1818181818F818F81818181818181818;
        8'hB6 : characterraster = 128'h36363636363636F63636363636363636;
        8'hB7 : characterraster = 128'h00000000000000FE3636363636363636;
        8'hB8 : characterraster = 128'h0000000000F818F81818181818181818;
        8'hB9 : characterraster = 128'h3636363636F606F63636363636363636;
        8'hBA : characterraster = 128'h36363636363636363636363636363636;
        8'hBB : characterraster = 128'h0000000000FE06F63636363636363636;
        8'hBC : characterraster = 128'h3636363636F606FE0000000000000000;
        8'hBD : characterraster = 128'h36363636363636FE0000000000000000;
        8'hBE : characterraster = 128'h1818181818F818F80000000000000000;
        8'hBF : characterraster = 128'h00000000000000F81818181818181818;
        8'hC0 : characterraster = 128'h181818181818181F0000000000000000;
        8'hC1 : characterraster = 128'h18181818181818FF0000000000000000;
        8'hC2 : characterraster = 128'h00000000000000FF1818181818181818;
        8'hC3 : characterraster = 128'h181818181818181F1818181818181818;
        8'hC4 : characterraster = 128'h00000000000000FF0000000000000000;
        8'hC5 : characterraster = 128'h18181818181818FF1818181818181818;
        8'hC6 : characterraster = 128'h18181818181F181F1818181818181818;
        8'hC7 : characterraster = 128'h36363636363636373636363636363636;
        8'hC8 : characterraster = 128'h363636363637303F0000000000000000;
        8'hC9 : characterraster = 128'h00000000003F30373636363636363636;
        8'hCA : characterraster = 128'h3636363636F700FF0000000000000000;
        8'hCB : characterraster = 128'h0000000000FF00F73636363636363636;
        8'hCC : characterraster = 128'h36363636363730373636363636363636;
        8'hCD : characterraster = 128'h0000000000FF00FF0000000000000000;
        8'hCE : characterraster = 128'h3636363636F700F73636363636363636;
        8'hCF : characterraster = 128'h1818181818FF00FF0000000000000000;
        8'hD0 : characterraster = 128'h36363636363636FF0000000000000000;
        8'hD1 : characterraster = 128'h0000000000FF00FF1818181818181818;
        8'hD2 : characterraster = 128'h00000000000000FF3636363636363636;
        8'hD3 : characterraster = 128'h363636363636363F0000000000000000;
        8'hD4 : characterraster = 128'h18181818181F181F0000000000000000;
        8'hD5 : characterraster = 128'h00000000001F181F1818181818181818;
        8'hD6 : characterraster = 128'h000000000000003F3636363636363636;
        8'hD7 : characterraster = 128'h36363636363636FF3636363636363636;
        8'hD8 : characterraster = 128'h1818181818FF18FF1818181818181818;
        8'hD9 : characterraster = 128'h18181818181818F80000000000000000;
        8'hDA : characterraster = 128'h000000000000001F1818181818181818;
        8'hDB : characterraster = 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
        8'hDC : characterraster = 128'h00000000000000FFFFFFFFFFFFFFFFFF;
        8'hDD : characterraster = 128'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0;
        8'hDE : characterraster = 128'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
        8'hDF : characterraster = 128'hFFFFFFFFFFFFFF000000000000000000;
        8'hE0 : characterraster = 128'h000000000076DCD8D8D8DC7600000000;
        8'hE1 : characterraster = 128'h000078CCCCCCD8CCC6C6C6CC00000000;
        8'hE2 : characterraster = 128'h0000FEC6C6C0C0C0C0C0C0C000000000;
        8'hE3 : characterraster = 128'h00000000FE6C6C6C6C6C6C6C00000000;
        8'hE4 : characterraster = 128'h000000FEC66030183060C6FE00000000;
        8'hE5 : characterraster = 128'h00000000007ED8D8D8D8D87000000000;
        8'hE6 : characterraster = 128'h0000000066666666667C6060C0000000;
        8'hE7 : characterraster = 128'h0000000076DC18181818181800000000;
        8'hE8 : characterraster = 128'h0000007E183C6666663C187E00000000;
        8'hE9 : characterraster = 128'h000000386CC6C6FEC6C66C3800000000;
        8'hEA : characterraster = 128'h0000386CC6C6C66C6C6C6CEE00000000;
        8'hEB : characterraster = 128'h00001E30180C3E666666663C00000000;
        8'hEC : characterraster = 128'h00000000007EDBDBDB7E000000000000;
        8'hED : characterraster = 128'h00000003067EDBDBF37E60C000000000;
        8'hEE : characterraster = 128'h00001C3060607C606060301C00000000;
        8'hEF : characterraster = 128'h0000007CC6C6C6C6C6C6C6C600000000;
        8'hF0 : characterraster = 128'h00000000FE0000FE0000FE0000000000;
        8'hF1 : characterraster = 128'h0000000018187E18180000FF00000000;
        8'hF2 : characterraster = 128'h00000030180C060C1830007E00000000;
        8'hF3 : characterraster = 128'h0000000C18306030180C007E00000000;
        8'hF4 : characterraster = 128'h00000E1B1B1818181818181818181818;
        8'hF5 : characterraster = 128'h1818181818181818D8D8D87000000000;
        8'hF6 : characterraster = 128'h000000001818007E0018180000000000;
        8'hF7 : characterraster = 128'h000000000076DC0076DC000000000000;
        8'hF8 : characterraster = 128'h00386C6C380000000000000000000000;
        8'hF9 : characterraster = 128'h00000000000000181800000000000000;
        8'hFA : characterraster = 128'h00000000000000001800000000000000;
        8'hFB : characterraster = 128'h000F0C0C0C0C0CEC6C6C3C1C00000000;
        8'hFC : characterraster = 128'h00D86C6C6C6C6C000000000000000000;
        8'hFD : characterraster = 128'h0070D83060C8F8000000000000000000;
        8'hFE : characterraster = 128'h000000007C7C7C7C7C7C7C0000000000;
        8'hFF : characterraster = 128'h00000000000000000000000000000000;
        default : characterraster = 0;
    endcase
end
endmodule
